module test(
    input logic CLK,
    input logic nRST,
    test_if.tuif tiif);
endmodule
